//test.sv
//description: test verilog files
//date: 2024-6-13

module new();

endmodule
